always @ (clk)
  begin
     ...     
  end // always @ (clk)
